**.subckt piezoresistor_tb
Xdut pres 0 vres 0 piezoresistor
Vres vres 0 1
Vpressure pres 0 0.9
**** begin user architecture code


.option savecurrents
.control
save all
dc vpressure 0.01 1.8 0.01 vres -2 2 1
write piezoresistor_tb.raw
plot all.Vres#branch
.endc


**** end user architecture code
**.ends

* expanding   symbol:  piezoresistor.sym # of pins=4
* sym_path: /home/cmaier/.xschem/sky130_TAC3/piezoresistor.sym
* sch_path: /home/cmaier/.xschem/sky130_TAC3/piezoresistor.sch
.subckt piezoresistor  pressure_pos pressure_neg resistor_pos resistor_neg
*.ipin pressure_pos
*.ipin pressure_neg
*.ipin resistor_pos
*.ipin resistor_neg
Broot sqrtp 0 V = sqrt(v(pressure_pos,pressure_neg))
Bres res 0 V = 106*(50/v(sqrtp)-1)*exp(-0.328*v(sqrtp))+15
Brvar resistor_pos resistor_neg I = V(resistor_pos,resistor_neg)/V(res)
.ends

** flattened .save nodes
.end
